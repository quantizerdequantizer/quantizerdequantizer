module Adder#(
   parameter WWIDTH  = 32,
   parameter WWIDTH_H  = 20
)(
   input  logic [0:0] clk,
   input  logic [WWIDTH-1:0] Mid,  
   input  logic [WWIDTH-1:0] ExtractedBits,
   output logic [WWIDTH-1:0] temp2,
   output logic              sign
);
logic [0:0] carry;
logic [WWIDTH-1:0] temp1;
logic [WWIDTH_H:0] temp1_H1;
logic [WWIDTH_H-1:0]  temp1_H2;
assign carry=temp1_H1[WWIDTH_H:WWIDTH_H];
always @(posedge clk) begin
	temp1_H1<= Mid[WWIDTH_H-1:0]+ExtractedBits[WWIDTH_H-1:0];
end
always @(posedge clk) begin
	temp1_H2<= Mid[WWIDTH-1:WWIDTH_H]+ExtractedBits[WWIDTH-1:WWIDTH_H]+carry;
end
assign temp1 = {temp1_H2,temp1_H1[WWIDTH_H-1:0]};
assign sign  = temp1[WWIDTH-1];
assign temp2 = sign ? temp1 : ~temp1 + 'h1; 
  
endmodule
